`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:25:50 04/12/2016 
// Design Name: 
// Module Name:    fourDigitDisplayTest 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module fourDigitDisplayTest(
    );

fourDigitDisplay display(clk_s, a_s, b_s, c_s, d_s, e_s, f_s, g_s, n3_s, n2_S, n1_s, n0_S);

endmodule
