`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:53:48 01/27/2015 
// Design Name: 
// Module Name:    votingtest 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
`timescale 1 ns/1 ns

module votingtest();

	reg s2, s1, s0, t, p;
	wire G;
	
	voting CompToTest(s2, s1, s0, t, p, G);
	
	initial begin
		// Test all possible input combinations
		s2 <= 0; s1 <= 0; s0 <= 0; t <= 0; p <= 0;    
		#10 s2 <= 0; s1 <= 0; s0 <= 0; t <= 0; p <= 1;      
		#10 s2 <= 0; s1 <= 0; s0 <= 0; t <= 1; p <= 0;      
		#10 s2 <= 0; s1 <= 0; s0 <= 0; t <= 1; p <= 1;     
		#10 s2 <= 0; s1 <= 0; s0 <= 1; t <= 0; p <= 0;        
		#10 s2 <= 0; s1 <= 0; s0 <= 1; t <= 0; p <= 1;        
		#10 s2 <= 0; s1 <= 0; s0 <= 1; t <= 1; p <= 0;         
		#10 s2 <= 0; s1 <= 0; s0 <= 1; t <= 1; p <= 1;       
		#10 s2 <= 0; s1 <= 1; s0 <= 0; t <= 0; p <= 0;          
		#10 s2 <= 0; s1 <= 1; s0 <= 0; t <= 0; p <= 1;      
		#10 s2 <= 0; s1 <= 1; s0 <= 0; t <= 1; p <= 0;     
		#10 s2 <= 0; s1 <= 1; s0 <= 0; t <= 1; p <= 1;        
		#10 s2 <= 0; s1 <= 1; s0 <= 1; t <= 0; p <= 0;       
		#10 s2 <= 0; s1 <= 1; s0 <= 1; t <= 0; p <= 1;        
		#10 s2 <= 0; s1 <= 1; s0 <= 1; t <= 1; p <= 0;       
		#10 s2 <= 0; s1 <= 1; s0 <= 1; t <= 1; p <= 1;        
		#10 s2 <= 1; s1 <= 0; s0 <= 0; t <= 0; p <= 0;        
		#10 s2 <= 1; s1 <= 0; s0 <= 0; t <= 0; p <= 1;        
		#10 s2 <= 1; s1 <= 0; s0 <= 0; t <= 1; p <= 0;        
		#10 s2 <= 1; s1 <= 0; s0 <= 0; t <= 1; p <= 1;         
		#10 s2 <= 1; s1 <= 0; s0 <= 1; t <= 0; p <= 0;     
		#10 s2 <= 1; s1 <= 0; s0 <= 1; t <= 0; p <= 1;        
		#10 s2 <= 1; s1 <= 0; s0 <= 1; t <= 1; p <= 0;     
		#10 s2 <= 1; s1 <= 0; s0 <= 1; t <= 1; p <= 1;        
		#10 s2 <= 1; s1 <= 1; s0 <= 0; t <= 0; p <= 0;         
		#10 s2 <= 1; s1 <= 1; s0 <= 0; t <= 0; p <= 1;         
		#10 s2 <= 1; s1 <= 1; s0 <= 0; t <= 1; p <= 0;        
		#10 s2 <= 1; s1 <= 1; s0 <= 0; t <= 1; p <= 1;        
		#10 s2 <= 1; s1 <= 1; s0 <= 1; t <= 0; p <= 0;        
		#10 s2 <= 1; s1 <= 1; s0 <= 1; t <= 0; p <= 1;     
		#10 s2 <= 1; s1 <= 1; s0 <= 1; t <= 1; p <= 0;       
		#10 s2 <= 1; s1 <= 1; s0 <= 1; t <= 1; p <= 1;
		
	end


endmodule


